// alu_opcodes.vh — ALU operation code definitions

`define ALU_ADD   5'd0
`define ALU_SUB   5'd1
`define ALU_AND   5'd2
`define ALU_OR    5'd3
`define ALU_XOR   5'd4
`define ALU_SLL   5'd5
`define ALU_SRL   5'd6
`define ALU_SRA   5'd7
`define ALU_SLT   5'd8
`define ALU_SLTU  5'd9
